* /home/shabbarvejlani/eSim-2.3/library/SubcircuitLibrary/epc_unit/epc_unit.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 08 Oct 2022 05:46:28 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
SC3  Net-_SC2-Pad1_ Net-_SC2-Pad2_ Net-_SC3-Pad3_ Net-_SC3-Pad4_ sky130_fd_pr__nfet_01v8		
SC4  Net-_SC3-Pad3_ Net-_SC4-Pad2_ Net-_SC3-Pad4_ Net-_SC3-Pad4_ sky130_fd_pr__nfet_01v8		
SC1  Net-_SC1-Pad1_ Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
SC2  Net-_SC2-Pad1_ Net-_SC2-Pad2_ Net-_SC1-Pad1_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
U1  Net-_SC1-Pad2_ Net-_SC2-Pad2_ Net-_SC4-Pad2_ Net-_SC3-Pad4_ Net-_SC1-Pad3_ Net-_SC2-Pad1_ PORT		

.end
